library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.all;

entity Data_memory is
    Port (
           clk : in std_logic;
           write : in std_logic;
           read : in std_logic;
           addr : in std_logic_vector (0 to 31);
           data_in : in std_logic_vector (0 to 31);
           
           data_out : out std_logic_vector (0 to 31)
           );
           end Data_memory;

architecture Behavioral of data_memory is

type MEM  is array (0 to 31) of std_logic_vector(0 to 31);

SIGNAL inst_mem: MEM :=(
"00000000000000000000000000000011","00000000000000000000000000000101",
"00000000000000000000000000000000","00000000000000000000000000000000",
"00000000000000000000000000000000","00000000000000000000000000000000",
"00000000000000000000000000000000","00000000000000000000000000000000",
"00000000000000000000000000000000","00000000000000000000000000000000",
"00000000000000000000000000000000","00000000000000000000000000000000",
"00000000000000000000000000000000","00000000000000000000000000000000",
"00000000000000000000000000000000","00000000000000000000000000000000",
"00000000000000000000000000000000","00000000000000000000000000000000",
"00000000000000000000000000000000","00000000000000000000000000000000",
"00000000000000000000000000000000","00000000000000000000000000000000",
"00000000000000000000000000000000","00000000000000000000000000000000",
"00000000000000000000000000000000","00000000000000000000000000000000",
"00000000000000000000000000000000","00000000000000000000000000000000",
"00000000000000000000000000000000","00000000000000000000000000000000",
"00000000000000000000000000000000","00000000000000000000000000000000"
);

begin 
    -- load
    data_out <= inst_mem(to_integer(unsigned(addr))) when read = '1';
    
    -- set
    inst_mem(to_integer(unsigned(addr))) <= data_in when write = '1' and rising_edge(clk); 

end Behavioral;